library IEEE;
use IEEE.STD_LOGIC_1164.all;
use ieee.numeric_std.all;


library work;
use work.trb_net_std.all;

entity delay_signal is
  generic(
    INPUT_WIDTH : integer;
    MAX_DEPTH   : integer
    );
  port(
    );
end entity;

architecture arch of delay_signal is

begin

end architecture;