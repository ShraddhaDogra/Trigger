library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.trb_net_std.all;
use work.trb_net_components.all;
use work.trb3_components.all;
use work.config.all;
use work.version.all;
use work.adc_package.all;

entity trb3sc_adc is
  port(
    --Clocks
    CLK_SUPPL_PCLK       : in    std_logic; --125 MHz for GbE
    CLK_CORE_PCLK        : in    std_logic; --Main Oscillator
    CLK_EXT_PLL_LEFT     : in    std_logic; --External Clock
    CLK_CORE_PLL_LEFT    : in    std_logic; --ADC Left 
    CLK_CORE_PLL_RIGHT   : in    std_logic; --ADC Right
    --Trigger
    TRIG_LEFT            : in    std_logic;  --left side trigger input from fan-out

    --Connection to AddOn               
    ADC1_CH              : in std_logic_vector(4 downto 0);
    ADC2_CH              : in std_logic_vector(4 downto 0);
    ADC3_CH              : in std_logic_vector(4 downto 0);
    ADC4_CH              : in std_logic_vector(4 downto 0);
    ADC5_CH              : in std_logic_vector(4 downto 0);
    ADC6_CH              : in std_logic_vector(4 downto 0);
    ADC7_CH              : in std_logic_vector(4 downto 0);
    ADC8_CH              : in std_logic_vector(4 downto 0);
    ADC9_CH              : in std_logic_vector(4 downto 0);
    ADC10_CH             : in std_logic_vector(4 downto 0);
    ADC11_CH             : in std_logic_vector(4 downto 0);
    ADC12_CH             : in std_logic_vector(4 downto 0);
    ADC_DCO              : in std_logic_vector(12 downto 1);

    SPI_ADC_SCK          : out std_logic;
    SPI_ADC_SDIO         : inout std_logic;
    
    LMK_CLK              : out std_logic;
    LMK_DATA             : out std_logic;
    LMK_LE_1             : out std_logic;
    LMK_LE_2             : out std_logic;
    
    P_CLOCK              : out std_logic;
    POWER_ENABLE         : out std_logic;
    
    FPGA_CS              : out std_logic_vector(1 downto 0);
    FPGA_SCK             : out std_logic_vector(1 downto 0);
    FPGA_SDI             : out std_logic_vector(1 downto 0);
    FPGA_SDO             : in  std_logic_vector(1 downto 0);
    
    
    --Additional IO
    HDR_IO               : inout std_logic_vector(10 downto 1);
    RJ_IO                : inout std_logic_vector( 3 downto 0);
    SPARE_IN             : in    std_logic_vector( 1 downto 0);  
    BACK_GPIO            : inout std_logic_vector( 3 downto 0);
    --LED
    LED_GREEN            : out   std_logic;
    LED_YELLOW           : out   std_logic;
    LED_ORANGE           : out   std_logic;
    LED_RED              : out   std_logic;
    LED_RJ_GREEN         : out   std_logic_vector( 1 downto 0);
    LED_RJ_RED           : out   std_logic_vector( 1 downto 0);
    LED_WHITE            : out   std_logic_vector( 1 downto 0);
    LED_SFP_GREEN        : out   std_logic_vector( 1 downto 0);
    LED_SFP_RED          : out   std_logic_vector( 1 downto 0);
    
    --SFP
    SFP_LOS              : in    std_logic_vector( 1 downto 0);
    SFP_MOD0             : in    std_logic_vector( 1 downto 0);  
    SFP_MOD1             : inout std_logic_vector( 1 downto 0) := (others => 'Z');
    SFP_MOD2             : inout std_logic_vector( 1 downto 0) := (others => 'Z');
    SFP_TX_DIS           : out   std_logic_vector( 1 downto 0) := (others => '0');  

    --Serdes switch
    PCSSW_ENSMB          : out   std_logic;
    PCSSW_EQ             : out   std_logic_vector( 3 downto 0);
    PCSSW_PE             : out   std_logic_vector( 3 downto 0);
    PCSSW                : out   std_logic_vector( 7 downto 0);
   
    --ADC
    ADC_CLK              : out   std_logic;
    ADC_CS               : out   std_logic;
    ADC_DIN              : out   std_logic;
    ADC_DOUT             : in    std_logic;

    --Flash, 1-wire, Reload
    FLASH_CLK            : out   std_logic;
    FLASH_CS             : out   std_logic;
    FLASH_IN             : out   std_logic;
    FLASH_OUT            : in    std_logic;
    PROGRAMN             : out   std_logic;
    ENPIRION_CLOCK       : out   std_logic;
    TEMPSENS             : inout std_logic;
    
    --Test Connectors
    TEST_LINE            : out std_logic_vector(15 downto 0)
    );
  attribute syn_useioff                  : boolean;
  --no IO-FF for LEDs relaxes timing constraints
  attribute syn_useioff of LED_GREEN     : signal is false;
  attribute syn_useioff of LED_ORANGE    : signal is false;
  attribute syn_useioff of LED_RED       : signal is false;
  attribute syn_useioff of LED_YELLOW    : signal is false;
  attribute syn_useioff of TEMPSENS      : signal is false;
  attribute syn_useioff of PROGRAMN      : signal is false;
  attribute syn_useioff of TRIG_LEFT     : signal is false;

  attribute syn_useioff of FLASH_CLK     : signal is true;
  attribute syn_useioff of FLASH_CS      : signal is true;
  attribute syn_useioff of FLASH_IN      : signal is true;
  attribute syn_useioff of FLASH_OUT     : signal is true;
  attribute syn_useioff of TEST_LINE     : signal is false;

  

end entity;


architecture trb3sc_adc_arch of trb3sc_adc is

  attribute syn_keep     : boolean;
  attribute syn_preserve : boolean;
  
  signal clk_sys, clk_full, clk_full_osc   : std_logic;
  signal GSR_N       : std_logic;
  signal reset_i     : std_logic;
  signal clear_i     : std_logic;
  
  signal time_counter      : unsigned(31 downto 0) := (others => '0');
  signal led               : std_logic_vector(1 downto 0);
  signal debug_clock_reset : std_logic_vector(31 downto 0);

  --Media Interface
  signal med2int           : med2int_array_t(0 to 0);
  signal int2med           : int2med_array_t(0 to 0);
  signal med_stat_debug    : std_logic_vector (1*64-1  downto 0);
  
  --READOUT
  signal readout_rx        : READOUT_RX;
  signal readout_tx        : readout_tx_array_t(0 to 11);

  signal ctrlbus_rx, bussci_rx, bustools_rx, bustc_rx, busadc_rx, bus_master_out  : CTRLBUS_RX;
  signal ctrlbus_tx, bussci_tx, bustools_tx, bustc_tx, busadc_tx, bus_master_in   : CTRLBUS_TX;
  
  signal common_stat_reg   : std_logic_vector(std_COMSTATREG*32-1 downto 0) := (others => '0');
  signal common_ctrl_reg   : std_logic_vector(std_COMCTRLREG*32-1 downto 0);
  
  signal sed_error_i       : std_logic;
  signal clock_select      : std_logic;
  signal bus_master_active : std_logic;
  
  signal spi_cs, spi_mosi, spi_miso, spi_clk : std_logic_vector(15 downto 0);

  signal timer    : TIMERS;
  signal lcd_data : std_logic_vector(511 downto 0);

  signal sfp_los_i, sfp_txdis_i, sfp_prsnt_i : std_logic;
  signal trig_gen_out_i : std_logic_vector(3 downto 0);

  signal adcspi_ctrl               : std_logic_vector(7 downto 0);

  signal s : std_logic_vector(3 downto 0);
attribute nopad : string;
attribute nopad of  s : signal is "true";  
  
begin
---------------------------------------------------------------------------
-- Clock & Reset Handling
---------------------------------------------------------------------------
THE_CLOCK_RESET :  entity work.clock_reset_handler
  port map(
    INT_CLK_IN      => CLK_CORE_PCLK,
    EXT_CLK_IN      => CLK_EXT_PLL_LEFT,
    NET_CLK_FULL_IN => med2int(0).clk_full,
    NET_CLK_HALF_IN => med2int(0).clk_half,
    RESET_FROM_NET  => med2int(0).stat_op(13),
    
    BUS_RX          => bustc_rx,
    BUS_TX          => bustc_tx,

    RESET_OUT       => reset_i,
    CLEAR_OUT       => clear_i,
    GSR_OUT         => GSR_N,
    
    FULL_CLK_OUT    => clk_full,
    SYS_CLK_OUT     => clk_sys,
    REF_CLK_OUT     => clk_full_osc,
    
    ENPIRION_CLOCK  => ENPIRION_CLOCK,    
    LED_RED_OUT     => LED_RJ_RED,
    LED_GREEN_OUT   => LED_RJ_GREEN,
    DEBUG_OUT       => debug_clock_reset
    );


---------------------------------------------------------------------------
-- TrbNet Uplink
---------------------------------------------------------------------------

  THE_MEDIA_INTERFACE : entity work.med_ecp3_sfp_sync
    generic map(
      SERDES_NUM    => SERDES_NUM,
      IS_SYNC_SLAVE => c_YES
      )
    port map(
      CLK_REF_FULL       => med2int(0).clk_full,
      CLK_INTERNAL_FULL  => clk_full_osc,
      SYSCLK        => clk_sys,
      RESET         => reset_i,
      CLEAR         => clear_i,
      --Internal Connection
      MEDIA_MED2INT => med2int(0),
      MEDIA_INT2MED => int2med(0),

      --Sync operation
      RX_DLM      => open,
      RX_DLM_WORD => open,
      TX_DLM      => open,
      TX_DLM_WORD => open,

      --SFP Connection
      SD_PRSNT_N_IN  => sfp_prsnt_i,
      SD_LOS_IN      => sfp_los_i,
      SD_TXDIS_OUT   => sfp_txdis_i,
      --Control Interface
      BUS_RX         => bussci_rx,
      BUS_TX         => bussci_tx,
      -- Status and control port
      STAT_DEBUG     => med_stat_debug(63 downto 0),
      CTRL_DEBUG     => open
      );


-- THE_MEDIA_INTERFACE_OLD : trb_net16_med_ecp3_sfp
--     generic map(
--       SERDES_NUM  => 0,        --number of serdes in quad
--       EXT_CLOCK   => c_NO,              --use internal clock
--       USE_200_MHZ => c_YES,             --run on 200 MHz clock
--       USE_125_MHZ => c_NO,
--       USE_CTC     => c_YES
--       )
--     port map(
--       CLK                => clk_full_osc,
--       SYSCLK             => clk_sys,
--       RESET              => reset_i,
--       CLEAR              => clear_i,
--       CLK_EN             => '1',
--       --Internal Connection
--       MED_DATA_IN        => int2med(0).data,
--       MED_PACKET_NUM_IN  => int2med(0).packet_num,
--       MED_DATAREADY_IN   => int2med(0).dataready,
--       MED_READ_OUT       => med2int(0).tx_read,
--       MED_DATA_OUT       => med2int(0).data,
--       MED_PACKET_NUM_OUT => med2int(0).packet_num,
--       MED_DATAREADY_OUT  => med2int(0).dataready,
--       MED_READ_IN        => '1',
--       REFCLK2CORE_OUT    => open,
--       --SFP Connection
--       SD_RXD_P_IN        => s(0),
--       SD_RXD_N_IN        => s(1),
--       SD_TXD_P_OUT       => s(2),
--       SD_TXD_N_OUT       => s(3),
--       SD_REFCLK_P_IN     => open,
--       SD_REFCLK_N_IN     => open,
--       SD_PRSNT_N_IN      => SFP_MOD0(0),
--       SD_LOS_IN          => SFP_LOS(0),
--       SD_TXDIS_OUT       => SFP_TX_DIS(0),
--       -- Status and control port
--       STAT_OP            => med2int(0).stat_op,
--       CTRL_OP            => int2med(0).ctrl_op,
--       STAT_DEBUG         => med_stat_debug(63 downto 0),
--       CTRL_DEBUG         => (others => '0')
--       );

  SFP_TX_DIS(0) <= '1';
  gen_sfp_con : if SERDES_NUM = 3 generate
    sfp_los_i   <= SFP_LOS(1);
    sfp_prsnt_i <= SFP_MOD0(1); 
    SFP_TX_DIS(1) <= sfp_txdis_i;
  end generate;  
  gen_bpl_con : if SERDES_NUM = 0 generate
    sfp_los_i   <= BACK_GPIO(1);
    sfp_prsnt_i <= BACK_GPIO(1); 
    BACK_GPIO(0) <= sfp_txdis_i;
  end generate;  
--   
---------------------------------------------------------------------------
-- Endpoint
---------------------------------------------------------------------------
THE_ENDPOINT : entity work.trb_net16_endpoint_hades_full_handler_record
  generic map (
    ADDRESS_MASK                 => x"FFFF",
    BROADCAST_BITMASK            => x"FF",
    REGIO_INIT_ENDPOINT_ID       => x"0001",
    TIMING_TRIGGER_RAW           => c_YES,
    --Configure data handler
      DATA_INTERFACE_NUMBER     => 12,
      DATA_BUFFER_DEPTH         => 10,
      DATA_BUFFER_WIDTH         => 32,
      DATA_BUFFER_FULL_THRESH   => 2**10-511,
      TRG_RELEASE_AFTER_DATA    => c_YES,
      HEADER_BUFFER_DEPTH       => 9,
      HEADER_BUFFER_FULL_THRESH => 2**9-16
      )
  port map(
    CLK                => clk_sys,
    RESET              => reset_i,
    CLK_EN             => '1',
    --  Media direction port
    MEDIA_MED2INT                => med2int(0),
    MEDIA_INT2MED                => int2med(0),
    --Timing trigger in
    TRG_TIMING_TRG_RECEIVED_IN   => TRIG_LEFT,
    READOUT_RX                   => readout_rx,
    READOUT_TX                   => readout_tx,

    --Slow Control Port
    REGIO_COMMON_STAT_REG_IN     => (others => '0'),  --0x00
    REGIO_COMMON_CTRL_REG_OUT    => common_ctrl_reg,  --0x20
    BUS_RX                       => ctrlbus_rx,
    BUS_TX                       => ctrlbus_tx,
    BUS_MASTER_IN                => bus_master_in,
    BUS_MASTER_OUT               => bus_master_out,
    BUS_MASTER_ACTIVE            => bus_master_active,   
    ONEWIRE_INOUT                => TEMPSENS,
    --Timing registers
    TIMERS_OUT                   => timer

    );

---------------------------------------------------------------------------
-- AddOn
---------------------------------------------------------------------------
gen_reallogic : if USE_DUMMY_READOUT = 0 generate
  THE_ADC : entity work.adc_handler
    generic map(
      IS_TRB3 = 0
      )
    port map(
      CLK        => clk_sys,
      CLK_ADCRAW => CLK_CORE_PCLK, --clk_full_osc,
      CLK_RAW_LEFT => CLK_CORE_PLL_LEFT,
      CLK_RAW_RIGHT=> CLK_CORE_PLL_RIGHT,

      ADCCLK_OUT => open, --P_CLOCK, 
      ADC_DATA( 4 downto  0)   => ADC1_CH,
      ADC_DATA( 9 downto  5)   => ADC2_CH,
      ADC_DATA(14 downto 10)   => ADC3_CH,
      ADC_DATA(19 downto 15)   => ADC4_CH,
      ADC_DATA(24 downto 20)   => ADC5_CH,
      ADC_DATA(29 downto 25)   => ADC6_CH,
      ADC_DATA(34 downto 30)   => ADC7_CH,
      ADC_DATA(39 downto 35)   => ADC8_CH,
      ADC_DATA(44 downto 40)   => ADC9_CH,
      ADC_DATA(49 downto 45)   => ADC10_CH,
      ADC_DATA(54 downto 50)   => ADC11_CH,
      ADC_DATA(59 downto 55)   => ADC12_CH,
      ADC_DCO     => ADC_DCO,
      TRIGGER_FLAG_OUT => trig_gen_out_i(0),
      
      TRIGGER_IN  => TRIG_LEFT,
      READOUT_RX  => readout_rx,
      READOUT_TX  => readout_tx,
      BUS_RX      => busadc_rx,
      BUS_TX      => busadc_tx,
      
      ADCSPI_CTRL => adcspi_ctrl
      );    
end generate;
    
gen_dummyreadout : if USE_DUMMY_READOUT = 1 generate
  THE_ADC : entity work.adc_slowcontrol_data_buffer
    port map(
      CLK        => clk_sys,
      CLK_ADCRAW => clk_full_osc,
      
      ADCCLK_OUT => open, --P_CLOCK,
      ADC_DATA( 4 downto  0)   => ADC1_CH,
      ADC_DATA( 9 downto  5)   => ADC2_CH,
      ADC_DATA(14 downto 10)   => ADC3_CH,
      ADC_DATA(19 downto 15)   => ADC4_CH,
      ADC_DATA(24 downto 20)   => ADC5_CH,
      ADC_DATA(29 downto 25)   => ADC6_CH,
      ADC_DATA(34 downto 30)   => ADC7_CH,
      ADC_DATA(39 downto 35)   => ADC8_CH,
      ADC_DATA(44 downto 40)   => ADC9_CH,
      ADC_DATA(49 downto 45)   => ADC10_CH,
      ADC_DATA(54 downto 50)   => ADC11_CH,
      ADC_DATA(59 downto 55)   => ADC12_CH,
      ADC_DCO     => ADC_DCO,
      
      ADC_CONTROL_OUT => adcspi_ctrl,
      
      BUS_RX      => busadc_rx,
      BUS_TX      => busadc_tx
      );
end generate;


  THE_ADC_REF : entity work.pll_in240_out40
    port map(
      CLK   => CLK_CORE_PCLK,
      CLKOP => P_CLOCK,
      LOCK  => open
      );
    
---------------------------------------------------------------------------
-- Bus Handler
---------------------------------------------------------------------------

  THE_BUS_HANDLER : entity work.trb_net16_regio_bus_handler_record
    generic map(
      PORT_NUMBER      => 4,
      PORT_ADDRESSES   => (0 => x"d000", 1 => x"b000", 2 => x"d300", 3 => x"a000", others => x"0000"),
      PORT_ADDR_MASK   => (0 => 12,      1 => 9,       2 => 1,       3 => 12,      others => 0),
      PORT_MASK_ENABLE => 1
      )
    port map(
      CLK   => clk_sys,
      RESET => reset_i,

      REGIO_RX  => ctrlbus_rx,
      REGIO_TX  => ctrlbus_tx,
      
      BUS_RX(0) => bustools_rx, --Flash, SPI, UART, ADC, SED
      BUS_RX(1) => bussci_rx,   --SCI Serdes
      BUS_RX(2) => bustc_rx,    --Clock switch
      BUS_RX(3) => busadc_rx,
      BUS_TX(0) => bustools_tx,
      BUS_TX(1) => bussci_tx,
      BUS_TX(2) => bustc_tx,
      BUS_TX(3) => busadc_tx,
      
      STAT_DEBUG => open
      );
      

---------------------------------------------------------------------------
-- Control Tools
---------------------------------------------------------------------------
  THE_TOOLS: entity work.trb3sc_tools 
    port map(
      CLK         => clk_sys,
      RESET       => reset_i,
      
      --Flash & Reload
      FLASH_CS    => FLASH_CS,
      FLASH_CLK   => FLASH_CLK,
      FLASH_IN    => FLASH_OUT,
      FLASH_OUT   => FLASH_IN,
      PROGRAMN    => PROGRAMN,
      REBOOT_IN   => common_ctrl_reg(15),
      --SPI
      SPI_CS_OUT  => spi_cs,  
      SPI_MOSI_OUT=> spi_mosi,
      SPI_MISO_IN => spi_miso,
      SPI_CLK_OUT => spi_clk,
      --Header
      HEADER_IO   => HDR_IO,
      --LCD
      LCD_DATA_IN => lcd_data,
      --ADC
      ADC_CS      => ADC_CS,
      ADC_MOSI    => ADC_DIN,
      ADC_MISO    => ADC_DOUT,
      ADC_CLK     => ADC_CLK,
      --SED
      SED_ERROR_OUT => sed_error_i,
      --Slowcontrol
      BUS_RX     => bustools_rx,
      BUS_TX     => bustools_tx,
      --Control master for default settings
      BUS_MASTER_IN  => bus_master_in,
      BUS_MASTER_OUT => bus_master_out,
      BUS_MASTER_ACTIVE => bus_master_active,      
      DEBUG_OUT  => open
      );

  -- the bits spi_CS (chip select) determines which SPI device is to be programmed
  -- it is already inverted, such that spi_CS=0xffff when nothing is to be programmed
  -- since the CS of the ADCs can only be controlled via the FPGA,
  -- we multiplex the SDI/O and SCK lines according to CS. This way we can control
  -- when which SPI device should be addressed via software

  FPGA_CS_mux: process (spi_cs(2 downto 0)) is
  begin  -- process FPGA_CS_mux
    case spi_cs(2 downto 0) is
      when b"110"  =>
        FPGA_CS <= b"00";
      when b"101"  =>
        FPGA_CS <= b"01";
      when b"011"  =>
        FPGA_CS <= b"10";        
      when others =>
        FPGA_CS <= b"11";
    end case;
  end process FPGA_CS_mux;
  
  FPGA_SCK(0) <= spi_clk(0)   when spi_cs(2 downto 0) /= b"111" else '1';
  FPGA_SDI(0) <= spi_mosi(0)  when spi_cs(2 downto 0) /= b"111" else '0';
  spi_miso(0) <= FPGA_SDO(0)  when spi_cs(2 downto 0) /= b"111" else '0';
  spi_miso(1) <= FPGA_SDO(0)  when spi_cs(2 downto 0) /= b"111" else '0';
  spi_miso(2) <= FPGA_SDO(0)  when spi_cs(2 downto 0) /= b"111" else '0';
  
  SPI_ADC_SCK         <= spi_clk(3)  when spi_cs(3) = '0' else adcspi_ctrl(4);
  SPI_ADC_SDIO        <= spi_mosi(3) when spi_cs(3) = '0' else adcspi_ctrl(5);
  FPGA_SCK(1)         <= '0'         when spi_cs(3) = '0' else adcspi_ctrl(6); --CSB
  
  LMK_CLK             <= spi_clk(4)  when spi_cs(5 downto 4) /= b"11" else '1' ;
  LMK_DATA            <= spi_mosi(4) when spi_cs(5 downto 4) /= b"11" else '0' ;
  LMK_LE_1            <= spi_cs(4); -- active low
  LMK_LE_2            <= spi_cs(5); -- active low
  
  POWER_ENABLE        <= adcspi_ctrl(0);

  
---------------------------------------------------------------------------
-- Switches
---------------------------------------------------------------------------
--Serdes Select
  PCSSW_ENSMB <= '0';
  PCSSW_EQ    <= x"0";
  PCSSW_PE    <= x"F";
  PCSSW       <= "01001110"; --SFP2 on B3, AddOn on D1

---------------------------------------------------------------------------
-- I/O
---------------------------------------------------------------------------

  RJ_IO(3 downto 2) <= trig_gen_out_i(1 downto 0);
  

  BACK_GPIO(1 downto 0)  <= (others => 'Z');
  BACK_GPIO(3 downto 2)  <= trig_gen_out_i(1 downto 0);
  
--   BACK_LVDS           <= (others => '0');
--   BACK_3V3            <= (others => 'Z');

  
---------------------------------------------------------------------------
-- LCD Data to display
---------------------------------------------------------------------------  
  lcd_data(15 downto 0)    <= timer.network_address;
  lcd_data(47 downto 16)   <= timer.microsecond;
  lcd_data(79 downto 48)   <= std_logic_vector(to_unsigned(VERSION_NUMBER_TIME,32));
  lcd_data(511 downto 80)  <= (others => '0');  
  
---------------------------------------------------------------------------
-- LED
---------------------------------------------------------------------------
  --LED are green, orange, red, yellow, white(2), rj_green(2), rj_red(2), sfp_green(2), sfp_red(2)
  LED_GREEN            <= debug_clock_reset(0);   
  LED_ORANGE           <= debug_clock_reset(1);
  LED_RED              <= not sed_error_i;
  LED_YELLOW           <= debug_clock_reset(2);
  LED_WHITE(0)         <= time_counter(26) and time_counter(19);  
  LED_WHITE(1)         <= time_counter(20);
  LED_SFP_GREEN        <= not med2int(0).stat_op(9) & '1';  --SFP Link Status
  LED_SFP_RED          <= not (med2int(0).stat_op(10) or med2int(0).stat_op(11)) & '1';  --SFP RX/TX

---------------------------------------------------------------------------
-- Test Circuits
---------------------------------------------------------------------------
  process begin
    wait until rising_edge(clk_sys);
    time_counter <= time_counter + 1; 
    if reset_i = '1' then
      time_counter <= (others => '0');
    end if;
  end process;  

  

end architecture;
