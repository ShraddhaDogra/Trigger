library ieee;
use ieee.std_logic_1164.all;
USE IEEE.numeric_std.ALL;
USE IEEE.std_logic_UNSIGNED.ALL;
library work;
use work.trb_net_std.all;

package trb_net_gbe_protocols is
	type hist_array is array (31 downto 0) of std_logic_vector(31 downto 0);

	--signal g_SIMULATE             : integer range 0 to 1 := 0;

	---- g_MY_IP is being set by DHCP Response Constructor
	--signal g_MY_IP                : std_logic_vector(31 downto 0);
	---- g_MY_MAC is being set by Main Controller
	--signal g_MY_MAC               : std_logic_vector(47 downto 0) := x"001122334455";

	constant c_MAX_FRAME_TYPES   : integer range 1 to 16 := 2;
	constant c_MAX_PROTOCOLS     : integer range 1 to 16 := 6; --5; --4; --5;
	constant c_MAX_IP_PROTOCOLS  : integer range 1 to 16 := 2;
	constant c_MAX_UDP_PROTOCOLS : integer range 1 to 16 := 4;

	type frame_types_a is array (c_MAX_FRAME_TYPES - 1 downto 0) of std_logic_vector(15 downto 0);
	constant FRAME_TYPES : frame_types_a := (x"0800", x"0806");
	-- IPv4, ARP

	type ip_protos_a is array (c_MAX_IP_PROTOCOLS - 1 downto 0) of std_logic_vector(7 downto 0);
	constant IP_PROTOCOLS : ip_protos_a := (x"11", x"01");
	-- UDP, ICMP

	-- this are the destination ports of the incoming packet
	type udp_protos_a is array (c_MAX_UDP_PROTOCOLS - 1 downto 0) of std_logic_vector(15 downto 0);
	constant UDP_PROTOCOLS : udp_protos_a := (x"0044", x"6590", x"7530", x"7531"); --x"6590", x"7530", x"7531"); --x"61a8", x"7530", x"7531");
	-- DHCP client, SCTRL, STATs

-- 	component trb_net16_gbe_response_constructor_Forward is
-- 	      port (
-- 		      CLK			: in	std_logic;  -- system clock
-- 		      RESET			: in	std_logic;
-- 		      
-- 	      -- INTERFACE	
-- 		      MY_MAC_IN                     : in  std_logic_vector(47 downto 0);
-- 		      MY_IP_IN                      : in  std_logic_vector(31 downto 0);
-- 		      PS_DATA_IN		: in	std_logic_vector(8 downto 0);
-- 		      PS_WR_EN_IN		: in	std_logic;
-- 		      PS_ACTIVATE_IN		: in	std_logic;
-- 		      PS_RESPONSE_READY_OUT	: out	std_logic;
-- 		      PS_BUSY_OUT		: out	std_logic;
-- 		      PS_SELECTED_IN		: in	std_logic;
-- 		      PS_SRC_MAC_ADDRESS_IN	: in	std_logic_vector(47 downto 0);
-- 		      PS_DEST_MAC_ADDRESS_IN  : in	std_logic_vector(47 downto 0);
-- 		      PS_SRC_IP_ADDRESS_IN	: in	std_logic_vector(31 downto 0);
-- 		      PS_DEST_IP_ADDRESS_IN	: in	std_logic_vector(31 downto 0);
-- 		      PS_SRC_UDP_PORT_IN	: in	std_logic_vector(15 downto 0);
-- 		      PS_DEST_UDP_PORT_IN	: in	std_logic_vector(15 downto 0);
-- 		      
-- 		      TC_RD_EN_IN		: in	std_logic;
-- 		      TC_DATA_OUT		: out	std_logic_vector(8 downto 0);
-- 		      TC_FRAME_SIZE_OUT	: out	std_logic_vector(15 downto 0);
-- 		      TC_FRAME_TYPE_OUT	: out	std_logic_vector(15 downto 0);
-- 		      TC_IP_PROTOCOL_OUT	: out	std_logic_vector(7 downto 0);	
-- 		      TC_DEST_MAC_OUT		: out	std_logic_vector(47 downto 0);
-- 		      TC_DEST_IP_OUT		: out	std_logic_vector(31 downto 0);
-- 		      TC_DEST_UDP_OUT		: out	std_logic_vector(15 downto 0);
-- 		      TC_SRC_MAC_OUT		: out	std_logic_vector(47 downto 0);
-- 		      TC_SRC_IP_OUT		: out	std_logic_vector(31 downto 0);
-- 		      TC_SRC_UDP_OUT		: out	std_logic_vector(15 downto 0);
-- 		      
-- 		      TC_BUSY_IN		: in	std_logic;
-- 			      
-- 		      RECEIVED_FRAMES_OUT	: out	std_logic_vector(15 downto 0);
-- 		      SENT_FRAMES_OUT		: out	std_logic_vector(15 downto 0);
-- 	      -- END OF INTERFACE
-- 
-- 		      FWD_DATA_IN		: in	std_logic_vector(7 downto 0);
-- 		      FWD_DATA_VALID_IN	: in	std_logic;
-- 		      FWD_SOP_IN		: in	std_logic;
-- 		      FWD_EOP_IN		: in	std_logic;
-- 		      FWD_READY_OUT		: out	std_logic;
-- 		      FWD_FULL_OUT		: out	std_logic;
-- 
-- 	      -- debug
-- 		      DEBUG_OUT		: out	std_logic_vector(31 downto 0)
-- 	      );
-- 	end component;

	component trb_net16_gbe_response_constructor_ARP is
		generic(STAT_ADDRESS_BASE : integer := 0
		);
		port(
			CLK                    : in  std_logic; -- system clock
			RESET                  : in  std_logic;

			-- INTERFACE	
			MY_MAC_IN              : in  std_logic_vector(47 downto 0);
			MY_IP_IN               : in  std_logic_vector(31 downto 0);
			PS_DATA_IN             : in  std_logic_vector(8 downto 0);
			PS_WR_EN_IN            : in  std_logic;
			PS_ACTIVATE_IN         : in  std_logic;
			PS_RESPONSE_READY_OUT  : out std_logic;
			PS_BUSY_OUT            : out std_logic;
			PS_SELECTED_IN         : in  std_logic;
			PS_SRC_MAC_ADDRESS_IN  : in  std_logic_vector(47 downto 0);
			PS_DEST_MAC_ADDRESS_IN : in  std_logic_vector(47 downto 0);
			PS_SRC_IP_ADDRESS_IN   : in  std_logic_vector(31 downto 0);
			PS_DEST_IP_ADDRESS_IN  : in  std_logic_vector(31 downto 0);
			PS_SRC_UDP_PORT_IN     : in  std_logic_vector(15 downto 0);
			PS_DEST_UDP_PORT_IN    : in  std_logic_vector(15 downto 0);
			TC_RD_EN_IN            : in  std_logic;
			TC_DATA_OUT            : out std_logic_vector(8 downto 0);
			TC_FRAME_SIZE_OUT      : out std_logic_vector(15 downto 0);
			TC_FRAME_TYPE_OUT      : out std_logic_vector(15 downto 0);
			TC_IP_PROTOCOL_OUT     : out std_logic_vector(7 downto 0);
			TC_IDENT_OUT           : out std_logic_vector(15 downto 0);
			TC_DEST_MAC_OUT        : out std_logic_vector(47 downto 0);
			TC_DEST_IP_OUT         : out std_logic_vector(31 downto 0);
			TC_DEST_UDP_OUT        : out std_logic_vector(15 downto 0);
			TC_SRC_MAC_OUT         : out std_logic_vector(47 downto 0);
			TC_SRC_IP_OUT          : out std_logic_vector(31 downto 0);
			TC_SRC_UDP_OUT         : out std_logic_vector(15 downto 0);
			STAT_DATA_OUT          : out std_logic_vector(31 downto 0);
			STAT_ADDR_OUT          : out std_logic_vector(7 downto 0);
			STAT_DATA_RDY_OUT      : out std_logic;
			STAT_DATA_ACK_IN       : in  std_logic;
			RECEIVED_FRAMES_OUT    : out std_logic_vector(15 downto 0);
			SENT_FRAMES_OUT        : out std_logic_vector(15 downto 0);
			-- END OF INTERFACE

			-- debug
			DEBUG_OUT              : out std_logic_vector(63 downto 0)
		);
	end component;

	component trb_net16_gbe_response_constructor_Test is
		port(
			CLK                    : in  std_logic; -- system clock
			RESET                  : in  std_logic;

			-- INTERFACE	
			MY_MAC_IN              : in  std_logic_vector(47 downto 0);
			MY_IP_IN               : in  std_logic_vector(31 downto 0);
			PS_DATA_IN             : in  std_logic_vector(8 downto 0);
			PS_WR_EN_IN            : in  std_logic;
			PS_ACTIVATE_IN         : in  std_logic;
			PS_RESPONSE_READY_OUT  : out std_logic;
			PS_BUSY_OUT            : out std_logic;
			PS_SELECTED_IN         : in  std_logic;
			PS_SRC_MAC_ADDRESS_IN  : in  std_logic_vector(47 downto 0);
			PS_DEST_MAC_ADDRESS_IN : in  std_logic_vector(47 downto 0);
			PS_SRC_IP_ADDRESS_IN   : in  std_logic_vector(31 downto 0);
			PS_DEST_IP_ADDRESS_IN  : in  std_logic_vector(31 downto 0);
			PS_SRC_UDP_PORT_IN     : in  std_logic_vector(15 downto 0);
			PS_DEST_UDP_PORT_IN    : in  std_logic_vector(15 downto 0);
			TC_WR_EN_OUT           : out std_logic;
			TC_DATA_OUT            : out std_logic_vector(8 downto 0);
			TC_FRAME_SIZE_OUT      : out std_logic_vector(15 downto 0);
			TC_FRAME_TYPE_OUT      : out std_logic_vector(15 downto 0);
			TC_IP_PROTOCOL_OUT     : out std_logic_vector(7 downto 0);
			TC_DEST_MAC_OUT        : out std_logic_vector(47 downto 0);
			TC_DEST_IP_OUT         : out std_logic_vector(31 downto 0);
			TC_DEST_UDP_OUT        : out std_logic_vector(15 downto 0);
			TC_SRC_MAC_OUT         : out std_logic_vector(47 downto 0);
			TC_SRC_IP_OUT          : out std_logic_vector(31 downto 0);
			TC_SRC_UDP_OUT         : out std_logic_vector(15 downto 0);
			TC_BUSY_IN             : in  std_logic;
			RECEIVED_FRAMES_OUT    : out std_logic_vector(15 downto 0);
			SENT_FRAMES_OUT        : out std_logic_vector(15 downto 0);
			-- END OF INTERFACE

			-- debug
			DEBUG_OUT              : out std_logic_vector(63 downto 0)
		);
	end component;

	component trb_net16_gbe_response_constructor_Trash is
		generic(STAT_ADDRESS_BASE : integer := 0
		);
		port(
			CLK                    : in  std_logic; -- system clock
			RESET                  : in  std_logic;

			-- INTERFACE
			MY_MAC_IN              : in  std_logic_vector(47 downto 0);
			MY_IP_IN               : in  std_logic_vector(31 downto 0);
			PS_DATA_IN             : in  std_logic_vector(8 downto 0);
			PS_WR_EN_IN            : in  std_logic;
			PS_ACTIVATE_IN         : in  std_logic;
			PS_RESPONSE_READY_OUT  : out std_logic;
			PS_BUSY_OUT            : out std_logic;
			PS_SELECTED_IN         : in  std_logic;
			PS_SRC_MAC_ADDRESS_IN  : in  std_logic_vector(47 downto 0);
			PS_DEST_MAC_ADDRESS_IN : in  std_logic_vector(47 downto 0);
			PS_SRC_IP_ADDRESS_IN   : in  std_logic_vector(31 downto 0);
			PS_DEST_IP_ADDRESS_IN  : in  std_logic_vector(31 downto 0);
			PS_SRC_UDP_PORT_IN     : in  std_logic_vector(15 downto 0);
			PS_DEST_UDP_PORT_IN    : in  std_logic_vector(15 downto 0);
			TC_RD_EN_IN            : in  std_logic;
			TC_DATA_OUT            : out std_logic_vector(8 downto 0);
			TC_FRAME_SIZE_OUT      : out std_logic_vector(15 downto 0);
			TC_SIZE_LEFT_OUT       : out std_logic_vector(15 downto 0);
			TC_FRAME_TYPE_OUT      : out std_logic_vector(15 downto 0);
			TC_IP_PROTOCOL_OUT     : out std_logic_vector(7 downto 0);
			TC_DEST_MAC_OUT        : out std_logic_vector(47 downto 0);
			TC_DEST_IP_OUT         : out std_logic_vector(31 downto 0);
			TC_DEST_UDP_OUT        : out std_logic_vector(15 downto 0);
			TC_SRC_MAC_OUT         : out std_logic_vector(47 downto 0);
			TC_SRC_IP_OUT          : out std_logic_vector(31 downto 0);
			TC_SRC_UDP_OUT         : out std_logic_vector(15 downto 0);
			TC_IDENT_OUT           : out std_logic_vector(15 downto 0);
			TC_IP_SIZE_OUT         : out std_logic_vector(15 downto 0);
			TC_UDP_SIZE_OUT        : out std_logic_vector(15 downto 0);
			TC_FLAGS_OFFSET_OUT    : out std_logic_vector(15 downto 0);
			TC_BUSY_IN             : in  std_logic;
			STAT_DATA_OUT          : out std_logic_vector(31 downto 0);
			STAT_ADDR_OUT          : out std_logic_vector(7 downto 0);
			STAT_DATA_RDY_OUT      : out std_logic;
			STAT_DATA_ACK_IN       : in  std_logic;
			RECEIVED_FRAMES_OUT    : out std_logic_vector(15 downto 0);
			SENT_FRAMES_OUT        : out std_logic_vector(15 downto 0);
			-- END OF INTERFACE

			-- debug
			DEBUG_OUT              : out std_logic_vector(63 downto 0)
		);
	end component;

	component trb_net16_gbe_response_constructor_DHCP is
		generic(
			STAT_ADDRESS_BASE : integer := 0;
			DO_SIMULATION     : integer := 0
		);
		port(
			CLK                    : in  std_logic; -- system clock
			RESET                  : in  std_logic;

			-- INTERFACE	
			MY_MAC_IN              : in  std_logic_vector(47 downto 0);
			MY_IP_IN               : in  std_logic_vector(31 downto 0);
			PS_DATA_IN             : in  std_logic_vector(8 downto 0);
			PS_WR_EN_IN            : in  std_logic;
			PS_ACTIVATE_IN         : in  std_logic;
			PS_RESPONSE_READY_OUT  : out std_logic;
			PS_BUSY_OUT            : out std_logic;
			PS_SELECTED_IN         : in  std_logic;
			PS_SRC_MAC_ADDRESS_IN  : in  std_logic_vector(47 downto 0);
			PS_DEST_MAC_ADDRESS_IN : in  std_logic_vector(47 downto 0);
			PS_SRC_IP_ADDRESS_IN   : in  std_logic_vector(31 downto 0);
			PS_DEST_IP_ADDRESS_IN  : in  std_logic_vector(31 downto 0);
			PS_SRC_UDP_PORT_IN     : in  std_logic_vector(15 downto 0);
			PS_DEST_UDP_PORT_IN    : in  std_logic_vector(15 downto 0);
			TC_RD_EN_IN            : in  std_logic;
			TC_DATA_OUT            : out std_logic_vector(8 downto 0);
			TC_FRAME_SIZE_OUT      : out std_logic_vector(15 downto 0);
			TC_FRAME_TYPE_OUT      : out std_logic_vector(15 downto 0);
			TC_IP_PROTOCOL_OUT     : out std_logic_vector(7 downto 0);
			TC_IDENT_OUT           : out std_logic_vector(15 downto 0);
			TC_DEST_MAC_OUT        : out std_logic_vector(47 downto 0);
			TC_DEST_IP_OUT         : out std_logic_vector(31 downto 0);
			TC_DEST_UDP_OUT        : out std_logic_vector(15 downto 0);
			TC_SRC_MAC_OUT         : out std_logic_vector(47 downto 0);
			TC_SRC_IP_OUT          : out std_logic_vector(31 downto 0);
			TC_SRC_UDP_OUT         : out std_logic_vector(15 downto 0);
			STAT_DATA_OUT          : out std_logic_vector(31 downto 0);
			STAT_ADDR_OUT          : out std_logic_vector(7 downto 0);
			STAT_DATA_RDY_OUT      : out std_logic;
			STAT_DATA_ACK_IN       : in  std_logic;
			RECEIVED_FRAMES_OUT    : out std_logic_vector(15 downto 0);
			SENT_FRAMES_OUT        : out std_logic_vector(15 downto 0);
			-- END OF INTERFACE

			MY_IP_OUT              : out std_logic_vector(31 downto 0);
			DHCP_START_IN          : in  std_logic;
			DHCP_DONE_OUT          : out std_logic;
			-- debug
			DEBUG_OUT              : out std_logic_vector(63 downto 0)
		);
	end component;

	component trb_net16_gbe_response_constructor_Ping is
		generic(STAT_ADDRESS_BASE : integer := 0
		);
		port(
			CLK                    : in  std_logic; -- system clock
			RESET                  : in  std_logic;

			-- INTERFACE	
			MY_MAC_IN              : in  std_logic_vector(47 downto 0);
			MY_IP_IN               : in  std_logic_vector(31 downto 0);
			PS_DATA_IN             : in  std_logic_vector(8 downto 0);
			PS_WR_EN_IN            : in  std_logic;
			PS_ACTIVATE_IN         : in  std_logic;
			PS_RESPONSE_READY_OUT  : out std_logic;
			PS_BUSY_OUT            : out std_logic;
			PS_SELECTED_IN         : in  std_logic;
			PS_SRC_MAC_ADDRESS_IN  : in  std_logic_vector(47 downto 0);
			PS_DEST_MAC_ADDRESS_IN : in  std_logic_vector(47 downto 0);
			PS_SRC_IP_ADDRESS_IN   : in  std_logic_vector(31 downto 0);
			PS_DEST_IP_ADDRESS_IN  : in  std_logic_vector(31 downto 0);
			PS_SRC_UDP_PORT_IN     : in  std_logic_vector(15 downto 0);
			PS_DEST_UDP_PORT_IN    : in  std_logic_vector(15 downto 0);
			TC_RD_EN_IN            : in  std_logic;
			TC_DATA_OUT            : out std_logic_vector(8 downto 0);
			TC_FRAME_SIZE_OUT      : out std_logic_vector(15 downto 0);
			TC_FRAME_TYPE_OUT      : out std_logic_vector(15 downto 0);
			TC_IP_PROTOCOL_OUT     : out std_logic_vector(7 downto 0);
			TC_IDENT_OUT           : out std_logic_vector(15 downto 0);
			TC_DEST_MAC_OUT        : out std_logic_vector(47 downto 0);
			TC_DEST_IP_OUT         : out std_logic_vector(31 downto 0);
			TC_DEST_UDP_OUT        : out std_logic_vector(15 downto 0);
			TC_SRC_MAC_OUT         : out std_logic_vector(47 downto 0);
			TC_SRC_IP_OUT          : out std_logic_vector(31 downto 0);
			TC_SRC_UDP_OUT         : out std_logic_vector(15 downto 0);
			STAT_DATA_OUT          : out std_logic_vector(31 downto 0);
			STAT_ADDR_OUT          : out std_logic_vector(7 downto 0);
			STAT_DATA_RDY_OUT      : out std_logic;
			STAT_DATA_ACK_IN       : in  std_logic;
			RECEIVED_FRAMES_OUT    : out std_logic_vector(15 downto 0);
			SENT_FRAMES_OUT        : out std_logic_vector(15 downto 0);
			-- END OF INTERFACE

			-- debug
			DEBUG_OUT              : out std_logic_vector(63 downto 0)
		);
	end component;
	
	component trb_net16_gbe_response_constructor_KillPing is
		generic(STAT_ADDRESS_BASE : integer := 0
		);
		port(
			CLK                    : in  std_logic; -- system clock
			RESET                  : in  std_logic;

			-- INTERFACE	
			MY_MAC_IN              : in  std_logic_vector(47 downto 0);
			MY_IP_IN               : in  std_logic_vector(31 downto 0);
			PS_DATA_IN             : in  std_logic_vector(8 downto 0);
			PS_WR_EN_IN            : in  std_logic;
			PS_ACTIVATE_IN         : in  std_logic;
			PS_RESPONSE_READY_OUT  : out std_logic;
			PS_BUSY_OUT            : out std_logic;
			PS_SELECTED_IN         : in  std_logic;
			PS_SRC_MAC_ADDRESS_IN  : in  std_logic_vector(47 downto 0);
			PS_DEST_MAC_ADDRESS_IN : in  std_logic_vector(47 downto 0);
			PS_SRC_IP_ADDRESS_IN   : in  std_logic_vector(31 downto 0);
			PS_DEST_IP_ADDRESS_IN  : in  std_logic_vector(31 downto 0);
			PS_SRC_UDP_PORT_IN     : in  std_logic_vector(15 downto 0);
			PS_DEST_UDP_PORT_IN    : in  std_logic_vector(15 downto 0);
			TC_RD_EN_IN            : in  std_logic;
			TC_DATA_OUT            : out std_logic_vector(8 downto 0);
			TC_FRAME_SIZE_OUT      : out std_logic_vector(15 downto 0);
			TC_FRAME_TYPE_OUT      : out std_logic_vector(15 downto 0);
			TC_IP_PROTOCOL_OUT     : out std_logic_vector(7 downto 0);
			TC_IDENT_OUT           : out std_logic_vector(15 downto 0);
			TC_DEST_MAC_OUT        : out std_logic_vector(47 downto 0);
			TC_DEST_IP_OUT         : out std_logic_vector(31 downto 0);
			TC_DEST_UDP_OUT        : out std_logic_vector(15 downto 0);
			TC_SRC_MAC_OUT         : out std_logic_vector(47 downto 0);
			TC_SRC_IP_OUT          : out std_logic_vector(31 downto 0);
			TC_SRC_UDP_OUT         : out std_logic_vector(15 downto 0);
			STAT_DATA_OUT          : out std_logic_vector(31 downto 0);
			STAT_ADDR_OUT          : out std_logic_vector(7 downto 0);
			STAT_DATA_RDY_OUT      : out std_logic;
			STAT_DATA_ACK_IN       : in  std_logic;
			RECEIVED_FRAMES_OUT    : out std_logic_vector(15 downto 0);
			SENT_FRAMES_OUT        : out std_logic_vector(15 downto 0);
			-- END OF INTERFACE
			
			MY_TRBNET_ADDRESS_IN : in std_logic_vector(15 downto 0);
			ISSUE_REBOOT_OUT : out std_logic;

			-- debug
			DEBUG_OUT              : out std_logic_vector(63 downto 0)
		);
	end component;

	component trb_net16_gbe_response_constructor_PseudoPing is
		generic(STAT_ADDRESS_BASE : integer := 0
		);
		port(
			CLK                    : in  std_logic; -- system clock
			RESET                  : in  std_logic;

			-- INTERFACE	
			MY_MAC_IN              : in  std_logic_vector(47 downto 0);
			MY_IP_IN               : in  std_logic_vector(31 downto 0);
			PS_DATA_IN             : in  std_logic_vector(8 downto 0);
			PS_WR_EN_IN            : in  std_logic;
			PS_ACTIVATE_IN         : in  std_logic;
			PS_RESPONSE_READY_OUT  : out std_logic;
			PS_BUSY_OUT            : out std_logic;
			PS_SELECTED_IN         : in  std_logic;
			PS_SRC_MAC_ADDRESS_IN  : in  std_logic_vector(47 downto 0);
			PS_DEST_MAC_ADDRESS_IN : in  std_logic_vector(47 downto 0);
			PS_SRC_IP_ADDRESS_IN   : in  std_logic_vector(31 downto 0);
			PS_DEST_IP_ADDRESS_IN  : in  std_logic_vector(31 downto 0);
			PS_SRC_UDP_PORT_IN     : in  std_logic_vector(15 downto 0);
			PS_DEST_UDP_PORT_IN    : in  std_logic_vector(15 downto 0);
			TC_RD_EN_IN            : in  std_logic;
			TC_DATA_OUT            : out std_logic_vector(8 downto 0);
			TC_FRAME_SIZE_OUT      : out std_logic_vector(15 downto 0);
			TC_FRAME_TYPE_OUT      : out std_logic_vector(15 downto 0);
			TC_IP_PROTOCOL_OUT     : out std_logic_vector(7 downto 0);
			TC_IDENT_OUT           : out std_logic_vector(15 downto 0);
			TC_DEST_MAC_OUT        : out std_logic_vector(47 downto 0);
			TC_DEST_IP_OUT         : out std_logic_vector(31 downto 0);
			TC_DEST_UDP_OUT        : out std_logic_vector(15 downto 0);
			TC_SRC_MAC_OUT         : out std_logic_vector(47 downto 0);
			TC_SRC_IP_OUT          : out std_logic_vector(31 downto 0);
			TC_SRC_UDP_OUT         : out std_logic_vector(15 downto 0);
			STAT_DATA_OUT          : out std_logic_vector(31 downto 0);
			STAT_ADDR_OUT          : out std_logic_vector(7 downto 0);
			STAT_DATA_RDY_OUT      : out std_logic;
			STAT_DATA_ACK_IN       : in  std_logic;
			RECEIVED_FRAMES_OUT    : out std_logic_vector(15 downto 0);
			SENT_FRAMES_OUT        : out std_logic_vector(15 downto 0);
			-- END OF INTERFACE

			-- debug
			DEBUG_OUT              : out std_logic_vector(63 downto 0)
		);
	end component;

	component trb_net16_gbe_response_constructor_Test1 is
		port(
			CLK                    : in  std_logic; -- system clock
			RESET                  : in  std_logic;

			-- INTERFACE	
			MY_MAC_IN              : in  std_logic_vector(47 downto 0);
			MY_IP_IN               : in  std_logic_vector(31 downto 0);
			PS_DATA_IN             : in  std_logic_vector(8 downto 0);
			PS_WR_EN_IN            : in  std_logic;
			PS_ACTIVATE_IN         : in  std_logic;
			PS_RESPONSE_READY_OUT  : out std_logic;
			PS_BUSY_OUT            : out std_logic;
			PS_SELECTED_IN         : in  std_logic;
			PS_SRC_MAC_ADDRESS_IN  : in  std_logic_vector(47 downto 0);
			PS_DEST_MAC_ADDRESS_IN : in  std_logic_vector(47 downto 0);
			PS_SRC_IP_ADDRESS_IN   : in  std_logic_vector(31 downto 0);
			PS_DEST_IP_ADDRESS_IN  : in  std_logic_vector(31 downto 0);
			PS_SRC_UDP_PORT_IN     : in  std_logic_vector(15 downto 0);
			PS_DEST_UDP_PORT_IN    : in  std_logic_vector(15 downto 0);
			TC_WR_EN_OUT           : out std_logic;
			TC_DATA_OUT            : out std_logic_vector(8 downto 0);
			TC_FRAME_SIZE_OUT      : out std_logic_vector(15 downto 0);
			TC_FRAME_TYPE_OUT      : out std_logic_vector(15 downto 0);
			TC_IP_PROTOCOL_OUT     : out std_logic_vector(7 downto 0);
			TC_DEST_MAC_OUT        : out std_logic_vector(47 downto 0);
			TC_DEST_IP_OUT         : out std_logic_vector(31 downto 0);
			TC_DEST_UDP_OUT        : out std_logic_vector(15 downto 0);
			TC_SRC_MAC_OUT         : out std_logic_vector(47 downto 0);
			TC_SRC_IP_OUT          : out std_logic_vector(31 downto 0);
			TC_SRC_UDP_OUT         : out std_logic_vector(15 downto 0);
			TC_BUSY_IN             : in  std_logic;
			RECEIVED_FRAMES_OUT    : out std_logic_vector(15 downto 0);
			SENT_FRAMES_OUT        : out std_logic_vector(15 downto 0);
			-- END OF INTERFACE

			-- debug
			DEBUG_OUT              : out std_logic_vector(63 downto 0)
		);
	end component;

	component trb_net16_gbe_response_constructor_SCTRL is
		generic(STAT_ADDRESS_BASE    : integer              := 0;
			    SLOWCTRL_BUFFER_SIZE : integer range 1 to 4 := 1
		);
		port(
			CLK                           : in  std_logic; -- system clock
			RESET                         : in  std_logic;

			-- INTERFACE	
			MY_MAC_IN                     : in  std_logic_vector(47 downto 0);
			MY_IP_IN                      : in  std_logic_vector(31 downto 0);
			PS_DATA_IN                    : in  std_logic_vector(8 downto 0);
			PS_WR_EN_IN                   : in  std_logic;
			PS_ACTIVATE_IN                : in  std_logic;
			PS_RESPONSE_READY_OUT         : out std_logic;
			PS_BUSY_OUT                   : out std_logic;
			PS_SELECTED_IN                : in  std_logic;
			PS_SRC_MAC_ADDRESS_IN         : in  std_logic_vector(47 downto 0);
			PS_DEST_MAC_ADDRESS_IN        : in  std_logic_vector(47 downto 0);
			PS_SRC_IP_ADDRESS_IN          : in  std_logic_vector(31 downto 0);
			PS_DEST_IP_ADDRESS_IN         : in  std_logic_vector(31 downto 0);
			PS_SRC_UDP_PORT_IN            : in  std_logic_vector(15 downto 0);
			PS_DEST_UDP_PORT_IN           : in  std_logic_vector(15 downto 0);
			TC_RD_EN_IN                   : in  std_logic;
			TC_DATA_OUT                   : out std_logic_vector(8 downto 0);
			TC_FRAME_SIZE_OUT             : out std_logic_vector(15 downto 0);
			TC_FRAME_TYPE_OUT             : out std_logic_vector(15 downto 0);
			TC_IP_PROTOCOL_OUT            : out std_logic_vector(7 downto 0);
			TC_IDENT_OUT                  : out std_logic_vector(15 downto 0);
			TC_DEST_MAC_OUT               : out std_logic_vector(47 downto 0);
			TC_DEST_IP_OUT                : out std_logic_vector(31 downto 0);
			TC_DEST_UDP_OUT               : out std_logic_vector(15 downto 0);
			TC_SRC_MAC_OUT                : out std_logic_vector(47 downto 0);
			TC_SRC_IP_OUT                 : out std_logic_vector(31 downto 0);
			TC_SRC_UDP_OUT                : out std_logic_vector(15 downto 0);
			STAT_DATA_OUT                 : out std_logic_vector(31 downto 0);
			STAT_ADDR_OUT                 : out std_logic_vector(7 downto 0);
			STAT_DATA_RDY_OUT             : out std_logic;
			STAT_DATA_ACK_IN              : in  std_logic;
			DEBUG_OUT                     : out std_logic_vector(63 downto 0);
			-- END OF INTERFACE

			-- protocol specific ports
			GSC_CLK_IN                    : in  std_logic;
			GSC_INIT_DATAREADY_OUT        : out std_logic;
			GSC_INIT_DATA_OUT             : out std_logic_vector(15 downto 0);
			GSC_INIT_PACKET_NUM_OUT       : out std_logic_vector(2 downto 0);
			GSC_INIT_READ_IN              : in  std_logic;
			GSC_REPLY_DATAREADY_IN        : in  std_logic;
			GSC_REPLY_DATA_IN             : in  std_logic_vector(15 downto 0);
			GSC_REPLY_PACKET_NUM_IN       : in  std_logic_vector(2 downto 0);
			GSC_REPLY_READ_OUT            : out std_logic;
			GSC_BUSY_IN                   : in  std_logic;
			MAKE_RESET_OUT                : out std_logic;
			CFG_ADDITIONAL_HDR_IN         : in  std_logic;
			CFG_MAX_REPLY_SIZE_IN         : in  std_logic_vector(31 downto 0);
			-- end of protocol specific ports

			MONITOR_SELECT_REC_OUT        : out std_logic_vector(31 downto 0);
			MONITOR_SELECT_REC_BYTES_OUT  : out std_logic_vector(31 downto 0);
			MONITOR_SELECT_SENT_BYTES_OUT : out std_logic_vector(31 downto 0);
			MONITOR_SELECT_SENT_OUT       : out std_logic_vector(31 downto 0);
			DATA_HIST_OUT                 : out hist_array
		);
	end component;

	component trb_net16_gbe_response_constructor_Stat is
		generic(STAT_ADDRESS_BASE : integer := 0
		);
		port(
			CLK                    : in  std_logic; -- system clock
			RESET                  : in  std_logic;

			-- INTERFACE	
			MY_MAC_IN              : in  std_logic_vector(47 downto 0);
			MY_IP_IN               : in  std_logic_vector(31 downto 0);
			PS_DATA_IN             : in  std_logic_vector(8 downto 0);
			PS_WR_EN_IN            : in  std_logic;
			PS_ACTIVATE_IN         : in  std_logic;
			PS_RESPONSE_READY_OUT  : out std_logic;
			PS_BUSY_OUT            : out std_logic;
			PS_SELECTED_IN         : in  std_logic;
			PS_SRC_MAC_ADDRESS_IN  : in  std_logic_vector(47 downto 0);
			PS_DEST_MAC_ADDRESS_IN : in  std_logic_vector(47 downto 0);
			PS_SRC_IP_ADDRESS_IN   : in  std_logic_vector(31 downto 0);
			PS_DEST_IP_ADDRESS_IN  : in  std_logic_vector(31 downto 0);
			PS_SRC_UDP_PORT_IN     : in  std_logic_vector(15 downto 0);
			PS_DEST_UDP_PORT_IN    : in  std_logic_vector(15 downto 0);
			TC_WR_EN_OUT           : out std_logic;
			TC_DATA_OUT            : out std_logic_vector(8 downto 0);
			TC_FRAME_SIZE_OUT      : out std_logic_vector(15 downto 0);
			TC_FRAME_TYPE_OUT      : out std_logic_vector(15 downto 0);
			TC_IP_PROTOCOL_OUT     : out std_logic_vector(7 downto 0);
			TC_IDENT_OUT           : out std_logic_vector(15 downto 0);
			TC_DEST_MAC_OUT        : out std_logic_vector(47 downto 0);
			TC_DEST_IP_OUT         : out std_logic_vector(31 downto 0);
			TC_DEST_UDP_OUT        : out std_logic_vector(15 downto 0);
			TC_SRC_MAC_OUT         : out std_logic_vector(47 downto 0);
			TC_SRC_IP_OUT          : out std_logic_vector(31 downto 0);
			TC_SRC_UDP_OUT         : out std_logic_vector(15 downto 0);
			TC_IP_SIZE_OUT         : out std_logic_vector(15 downto 0);
			TC_UDP_SIZE_OUT        : out std_logic_vector(15 downto 0);
			TC_FLAGS_OFFSET_OUT    : out std_logic_vector(15 downto 0);
			TC_BUSY_IN             : in  std_logic;
			STAT_DATA_OUT          : out std_logic_vector(31 downto 0);
			STAT_ADDR_OUT          : out std_logic_vector(7 downto 0);
			STAT_DATA_RDY_OUT      : out std_logic;
			STAT_DATA_ACK_IN       : in  std_logic;
			RECEIVED_FRAMES_OUT    : out std_logic_vector(15 downto 0);
			SENT_FRAMES_OUT        : out std_logic_vector(15 downto 0);
			-- END OF INTERFACE

			STAT_DATA_IN           : in  std_logic_vector((c_MAX_PROTOCOLS + 1) * 32 - 1 downto 0);
			STAT_ADDR_IN           : in  std_logic_vector((c_MAX_PROTOCOLS + 1) * 8 - 1 downto 0);
			STAT_DATA_RDY_IN       : in  std_logic_vector((c_MAX_PROTOCOLS + 1) - 1 downto 0);
			STAT_DATA_ACK_OUT      : out std_logic_vector((c_MAX_PROTOCOLS + 1) - 1 downto 0);

			-- debug
			DEBUG_OUT              : out std_logic_vector(63 downto 0)
		);
	end component;

	component trb_net16_gbe_response_constructor_TrbNetData is
		generic(
			RX_PATH_ENABLE      : integer range 0 to 1 := 1;
			DO_SIMULATION       : integer range 0 to 1 := 0;
			READOUT_BUFFER_SIZE : integer range 1 to 4 := 1
		);
		port(
			CLK                           : in  std_logic; -- system clock
			RESET                         : in  std_logic;

			-- INTERFACE	
			MY_MAC_IN                     : in  std_logic_vector(47 downto 0);
			MY_IP_IN                      : in  std_logic_vector(31 downto 0);
			PS_DATA_IN                    : in  std_logic_vector(8 downto 0);
			PS_WR_EN_IN                   : in  std_logic;
			PS_ACTIVATE_IN                : in  std_logic;
			PS_RESPONSE_READY_OUT         : out std_logic;
			PS_BUSY_OUT                   : out std_logic;
			PS_SELECTED_IN                : in  std_logic;
			PS_SRC_MAC_ADDRESS_IN         : in  std_logic_vector(47 downto 0);
			PS_DEST_MAC_ADDRESS_IN        : in  std_logic_vector(47 downto 0);
			PS_SRC_IP_ADDRESS_IN          : in  std_logic_vector(31 downto 0);
			PS_DEST_IP_ADDRESS_IN         : in  std_logic_vector(31 downto 0);
			PS_SRC_UDP_PORT_IN            : in  std_logic_vector(15 downto 0);
			PS_DEST_UDP_PORT_IN           : in  std_logic_vector(15 downto 0);
			TC_RD_EN_IN                   : in  std_logic;
			TC_DATA_OUT                   : out std_logic_vector(8 downto 0);
			TC_FRAME_SIZE_OUT             : out std_logic_vector(15 downto 0);
			TC_FRAME_TYPE_OUT             : out std_logic_vector(15 downto 0);
			TC_IP_PROTOCOL_OUT            : out std_logic_vector(7 downto 0);
			TC_IDENT_OUT                  : out std_logic_vector(15 downto 0);
			TC_DEST_MAC_OUT               : out std_logic_vector(47 downto 0);
			TC_DEST_IP_OUT                : out std_logic_vector(31 downto 0);
			TC_DEST_UDP_OUT               : out std_logic_vector(15 downto 0);
			TC_SRC_MAC_OUT                : out std_logic_vector(47 downto 0);
			TC_SRC_IP_OUT                 : out std_logic_vector(31 downto 0);
			TC_SRC_UDP_OUT                : out std_logic_vector(15 downto 0);
			STAT_DATA_OUT                 : out std_logic_vector(31 downto 0);
			STAT_ADDR_OUT                 : out std_logic_vector(7 downto 0);
			STAT_DATA_RDY_OUT             : out std_logic;
			STAT_DATA_ACK_IN              : in  std_logic;
			DEBUG_OUT                     : out std_logic_vector(63 downto 0);

			-- END OF INTERFACE

			-- CTS interface
			CTS_NUMBER_IN                 : in  std_logic_vector(15 downto 0);
			CTS_CODE_IN                   : in  std_logic_vector(7 downto 0);
			CTS_INFORMATION_IN            : in  std_logic_vector(7 downto 0);
			CTS_READOUT_TYPE_IN           : in  std_logic_vector(3 downto 0);
			CTS_START_READOUT_IN          : in  std_logic;
			CTS_DATA_OUT                  : out std_logic_vector(31 downto 0);
			CTS_DATAREADY_OUT             : out std_logic;
			CTS_READOUT_FINISHED_OUT      : out std_logic;
			CTS_READ_IN                   : in  std_logic;
			CTS_LENGTH_OUT                : out std_logic_vector(15 downto 0);
			CTS_ERROR_PATTERN_OUT         : out std_logic_vector(31 downto 0);
			-- Data payload interface
			FEE_DATA_IN                   : in  std_logic_vector(15 downto 0);
			FEE_DATAREADY_IN              : in  std_logic;
			FEE_READ_OUT                  : out std_logic;
			FEE_STATUS_BITS_IN            : in  std_logic_vector(31 downto 0);
			FEE_BUSY_IN                   : in  std_logic;
			-- ip configurator
			SLV_ADDR_IN                   : in  std_logic_vector(7 downto 0);
			SLV_READ_IN                   : in  std_logic;
			SLV_WRITE_IN                  : in  std_logic;
			SLV_BUSY_OUT                  : out std_logic;
			SLV_ACK_OUT                   : out std_logic;
			SLV_DATA_IN                   : in  std_logic_vector(31 downto 0);
			SLV_DATA_OUT                  : out std_logic_vector(31 downto 0);
			CFG_GBE_ENABLE_IN             : in  std_logic;
			CFG_IPU_ENABLE_IN             : in  std_logic;
			CFG_MULT_ENABLE_IN            : in  std_logic;
			CFG_SUBEVENT_ID_IN            : in  std_logic_vector(31 downto 0);
			CFG_SUBEVENT_DEC_IN           : in  std_logic_vector(31 downto 0);
			CFG_QUEUE_DEC_IN              : in  std_logic_vector(31 downto 0);
			CFG_READOUT_CTR_IN            : in  std_logic_vector(23 downto 0);
			CFG_READOUT_CTR_VALID_IN      : in  std_logic;
			CFG_INSERT_TTYPE_IN           : in  std_logic;
			CFG_MAX_SUB_IN                : in  std_logic_vector(15 downto 0);
			CFG_MAX_QUEUE_IN              : in  std_logic_vector(15 downto 0);
			CFG_MAX_SUBS_IN_QUEUE_IN      : in  std_logic_vector(15 downto 0);
			CFG_MAX_SINGLE_SUB_IN         : in  std_logic_vector(15 downto 0);
			CFG_AUTO_THROTTLE_IN          : in  std_logic;
			CFG_THROTTLE_PAUSE_IN         : in  std_logic_vector(15 downto 0);
			MONITOR_SELECT_REC_OUT        : out std_logic_vector(31 downto 0);
			MONITOR_SELECT_REC_BYTES_OUT  : out std_logic_vector(31 downto 0);
			MONITOR_SELECT_SENT_BYTES_OUT : out std_logic_vector(31 downto 0);
			MONITOR_SELECT_SENT_OUT       : out std_logic_vector(31 downto 0);
			MONITOR_SELECT_DROP_IN_OUT    : out std_logic_vector(31 downto 0);
			MONITOR_SELECT_DROP_OUT_OUT   : out std_logic_vector(31 downto 0);
			DATA_HIST_OUT                 : out hist_array
		);
	end component;

end package;
